�� sr Student'{@��OX I ageL 	firstNamet Ljava/lang/String;L lastNameq ~ xp   t Ivant Ivanov